x"018a",
x"0188",
x"048b",
x"048c",
x"008e",
x"010e",
x"090b",
x"048c",
x"048d",
x"090d",
x"0009",
