x"008e",
x"010e",
x"018e",
x"020e",
x"0e90",
x"8611",
x"9712",
x"9e13",
x"4154",
x"ffff",
x"4511",